typedef class nathiya;
  class nalinaa;
    nathiya y;
  endclass
  class nathiya;
    nalinaa l;
  endclass
  module typedef_class;
    initial
      begin
      
    $display("inside module");
    end
  endmodule
