module assosiative_array;
  int array1[int];
  int array2[string];
  int array3[string];
  initial
    begin
      array1='{1:22,6:34};
      array2='{"rose":100,"oey":200};
      array3='{"apple":"orange","pears":"44"};
  $display("array1=%p",array1);
      $display("array2=%p",array2);
      $display("array3=%p",array3);
  end
endmodule
